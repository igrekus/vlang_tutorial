module main

import cmod

fn main() {
	println('hi')
	cmod.hello_from_cmod()
	cmod.hello_from_c()
}
