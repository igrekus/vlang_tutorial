module mymod

pub fn impl_fn() {
	println('impl fn')
}
