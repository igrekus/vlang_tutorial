module tests_example

fn test_hello() {
	assert hello() == 'hello world'
}
